module SIPO_CB(CLOCK_CB, EN_CB, RES_CB, DAT_IN_CB, DAT_OUT_CB);

input CLOCK_CB, EN_CB, RES_CB, DAT_IN_CB;
output reg[111:0]DAT_OUT_CB;

always@(posedge CLOCK_CB)
if(~RES_CB)
begin
if(EN_CB)
begin
  DAT_OUT_CB[111]<=DAT_IN_CB;   
  DAT_OUT_CB[110]<=DAT_OUT_CB[111];
  DAT_OUT_CB[109]<=DAT_OUT_CB[110];
  DAT_OUT_CB[108]<=DAT_OUT_CB[109];
  DAT_OUT_CB[107]<=DAT_OUT_CB[108];
  DAT_OUT_CB[106]<=DAT_OUT_CB[107];
  DAT_OUT_CB[105]<=DAT_OUT_CB[106];
  DAT_OUT_CB[104]<=DAT_OUT_CB[105];
  DAT_OUT_CB[103]<=DAT_OUT_CB[104];
  DAT_OUT_CB[102]<=DAT_OUT_CB[103];
  DAT_OUT_CB[101]<=DAT_OUT_CB[102];
  DAT_OUT_CB[100]<=DAT_OUT_CB[101];
  DAT_OUT_CB[99]<=DAT_OUT_CB[100];
  DAT_OUT_CB[98]<=DAT_OUT_CB[99];
  DAT_OUT_CB[97]<=DAT_OUT_CB[98];
  DAT_OUT_CB[96]<=DAT_OUT_CB[97];
  DAT_OUT_CB[95]<=DAT_OUT_CB[96];
  DAT_OUT_CB[94]<=DAT_OUT_CB[95];
  DAT_OUT_CB[93]<=DAT_OUT_CB[94];
  DAT_OUT_CB[92]<=DAT_OUT_CB[93];
  DAT_OUT_CB[91]<=DAT_OUT_CB[92];
  DAT_OUT_CB[90]<=DAT_OUT_CB[91];
  DAT_OUT_CB[89]<=DAT_OUT_CB[90];
  DAT_OUT_CB[88]<=DAT_OUT_CB[89];
  DAT_OUT_CB[87]<=DAT_OUT_CB[88];
  DAT_OUT_CB[86]<=DAT_OUT_CB[87];
  DAT_OUT_CB[85]<=DAT_OUT_CB[86];
  DAT_OUT_CB[84]<=DAT_OUT_CB[85];
  DAT_OUT_CB[83]<=DAT_OUT_CB[84];
  DAT_OUT_CB[82]<=DAT_OUT_CB[83];
  DAT_OUT_CB[81]<=DAT_OUT_CB[82];
  DAT_OUT_CB[80]<=DAT_OUT_CB[81];
  DAT_OUT_CB[79]<=DAT_OUT_CB[80];
  DAT_OUT_CB[78]<=DAT_OUT_CB[79];
  DAT_OUT_CB[77]<=DAT_OUT_CB[78];
  DAT_OUT_CB[76]<=DAT_OUT_CB[77];
  DAT_OUT_CB[75]<=DAT_OUT_CB[76];
  DAT_OUT_CB[74]<=DAT_OUT_CB[75];
  DAT_OUT_CB[73]<=DAT_OUT_CB[74];
  DAT_OUT_CB[72]<=DAT_OUT_CB[73]; 
  DAT_OUT_CB[71]<=DAT_OUT_CB[72];
  DAT_OUT_CB[70]<=DAT_OUT_CB[71];
  DAT_OUT_CB[69]<=DAT_OUT_CB[70];
  DAT_OUT_CB[68]<=DAT_OUT_CB[69];
  DAT_OUT_CB[67]<=DAT_OUT_CB[68];
  DAT_OUT_CB[66]<=DAT_OUT_CB[67];
  DAT_OUT_CB[65]<=DAT_OUT_CB[66];
  DAT_OUT_CB[64]<=DAT_OUT_CB[65];
  DAT_OUT_CB[63]<=DAT_OUT_CB[64];
  DAT_OUT_CB[62]<=DAT_OUT_CB[63];
  DAT_OUT_CB[61]<=DAT_OUT_CB[62];
  DAT_OUT_CB[60]<=DAT_OUT_CB[61];
  DAT_OUT_CB[59]<=DAT_OUT_CB[60];
  DAT_OUT_CB[58]<=DAT_OUT_CB[59];
  DAT_OUT_CB[57]<=DAT_OUT_CB[58];
  DAT_OUT_CB[56]<=DAT_OUT_CB[57];
  DAT_OUT_CB[55]<=DAT_OUT_CB[56];
  DAT_OUT_CB[54]<=DAT_OUT_CB[55];
  DAT_OUT_CB[53]<=DAT_OUT_CB[54];
  DAT_OUT_CB[52]<=DAT_OUT_CB[53];
  DAT_OUT_CB[51]<=DAT_OUT_CB[52];
  DAT_OUT_CB[50]<=DAT_OUT_CB[51];
  DAT_OUT_CB[49]<=DAT_OUT_CB[50];
  DAT_OUT_CB[48]<=DAT_OUT_CB[49];
  DAT_OUT_CB[47]<=DAT_OUT_CB[48];
  DAT_OUT_CB[46]<=DAT_OUT_CB[47];
  DAT_OUT_CB[45]<=DAT_OUT_CB[46];
  DAT_OUT_CB[44]<=DAT_OUT_CB[45];
  DAT_OUT_CB[43]<=DAT_OUT_CB[44];
  DAT_OUT_CB[42]<=DAT_OUT_CB[43];
  DAT_OUT_CB[41]<=DAT_OUT_CB[42];
  DAT_OUT_CB[40]<=DAT_OUT_CB[41];
  DAT_OUT_CB[39]<=DAT_OUT_CB[40];
  DAT_OUT_CB[38]<=DAT_OUT_CB[39];
  DAT_OUT_CB[37]<=DAT_OUT_CB[38];
  DAT_OUT_CB[36]<=DAT_OUT_CB[37];
  DAT_OUT_CB[35]<=DAT_OUT_CB[36];
  DAT_OUT_CB[34]<=DAT_OUT_CB[35];
  DAT_OUT_CB[33]<=DAT_OUT_CB[34];
  DAT_OUT_CB[32]<=DAT_OUT_CB[33];
  DAT_OUT_CB[31]<=DAT_OUT_CB[32];
  DAT_OUT_CB[30]<=DAT_OUT_CB[31];
  DAT_OUT_CB[29]<=DAT_OUT_CB[30];
  DAT_OUT_CB[28]<=DAT_OUT_CB[29];
  DAT_OUT_CB[27]<=DAT_OUT_CB[28];
  DAT_OUT_CB[26]<=DAT_OUT_CB[27];
  DAT_OUT_CB[25]<=DAT_OUT_CB[26];
  DAT_OUT_CB[24]<=DAT_OUT_CB[25];
  DAT_OUT_CB[23]<=DAT_OUT_CB[24];
  DAT_OUT_CB[22]<=DAT_OUT_CB[23];
  DAT_OUT_CB[21]<=DAT_OUT_CB[22];
  DAT_OUT_CB[20]<=DAT_OUT_CB[21];
  DAT_OUT_CB[19]<=DAT_OUT_CB[20];
  DAT_OUT_CB[18]<=DAT_OUT_CB[19];
  DAT_OUT_CB[17]<=DAT_OUT_CB[18];
  DAT_OUT_CB[16]<=DAT_OUT_CB[17];
  DAT_OUT_CB[15]<=DAT_OUT_CB[16];
  DAT_OUT_CB[14]<=DAT_OUT_CB[15];
  DAT_OUT_CB[13]<=DAT_OUT_CB[14];
  DAT_OUT_CB[12]<=DAT_OUT_CB[13];
  DAT_OUT_CB[11]<=DAT_OUT_CB[12];
  DAT_OUT_CB[10]<=DAT_OUT_CB[11];
  DAT_OUT_CB[9]<=DAT_OUT_CB[10];
  DAT_OUT_CB[8]<=DAT_OUT_CB[9];
  DAT_OUT_CB[7]<=DAT_OUT_CB[8];
  DAT_OUT_CB[6]<=DAT_OUT_CB[7];
  DAT_OUT_CB[5]<=DAT_OUT_CB[6];
  DAT_OUT_CB[4]<=DAT_OUT_CB[5];
  DAT_OUT_CB[3]<=DAT_OUT_CB[4];
  DAT_OUT_CB[2]<=DAT_OUT_CB[3];
  DAT_OUT_CB[1]<=DAT_OUT_CB[2];
  DAT_OUT_CB[0]<=DAT_OUT_CB[1];
end
else
begin
  DAT_OUT_CB = DAT_OUT_CB;
end
end
else
begin
  DAT_OUT_CB = 1'b0;
end
endmodule
